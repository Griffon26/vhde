entity used_entity is
  port (
    myport1: in sometype;
    myport2: inout sometype
  );
end used_entity;

architecture used_arch of used_entity is


begin
end;
